module tb_alu();

endmodule
