module tb_adder();

endmodule
